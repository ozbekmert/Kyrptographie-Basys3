LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

LIBRARY UNISIM;
USE UNISIM.VCOMPONENTS.ALL;


ENTITY RegisterSerPar is
	GENERIC ( SIZE_SER	: POSITIVE := 1;
				 SIZE_PAR	: POSITIVE := 8);
	PORT ( CLK 	: IN  STD_LOGIC;
		   RST	: IN  STD_LOGIC;
           EN 	: IN  STD_LOGIC;
           SEL 	: IN  STD_LOGIC;
           DS 	: IN  STD_LOGIC_VECTOR((SIZE_SER - 1) DOWNTO 0);
           DP 	: IN  STD_LOGIC_VECTOR((SIZE_PAR - 1) DOWNTO 0);
           QS 	: OUT STD_LOGIC_VECTOR((SIZE_SER - 1) DOWNTO 0);
           QP 	: OUT STD_LOGIC_VECTOR((SIZE_PAR - 1) DOWNTO 0));
END RegisterSerPar;



ARCHITECTURE Mixed OF RegisterSerPar IS

    SIGNAL DP_INTERN, QP_INTERN : STD_LOGIC_VECTOR ((SIZE_PAR - 1) DOWNTO 0);

BEGIN

	DP_INTERN <= QP_INTERN ((SIZE_PAR - SIZE_SER - 1) DOWNTO 0) & DS WHEN (SEL = '0') ELSE DP;

	GEN :
	FOR I IN 0 TO (SIZE_PAR - 1) GENERATE
		FF : FDRE
		PORT MAP (
			C 	=> CLK,
			R	=> RST,
			CE	=> EN,
			D	=> DP_INTERN(I),
			Q	=> QP_INTERN(I)
		);
	END GENERATE;

	QS <= QP_INTERN((SIZE_PAR - 1) DOWNTO (SIZE_PAR - SIZE_SER));
	QP <= QP_INTERN;
	
END Mixed;

